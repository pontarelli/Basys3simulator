`timescale 1ns / 1ps

module ball_rom(
    input [2:0] addr,   // 3-bit address
    output reg [7:0] data   // 8-bit data
    );
    
    always @*
        case(addr)
            3'b000 :    data = 8'b00100100; //   ****  
            3'b001 :    data = 8'b01100110; //  ******
            3'b010 :    data = 8'b11100111; // ********
            3'b011 :    data = 8'b00000000; // ********
            3'b100 :    data = 8'b00000000; // ********
            3'b101 :    data = 8'b11100111; // ********
            3'b110 :    data = 8'b01100110; //  ******
            3'b111 :    data = 8'b00100100; //   ****
        endcase
    
endmodule

module ball_rom4(
    input [3:0] addr,   // 4-bit address
    output reg [15:0] data   // 16-bit data
    );
    
    always @*
        case(addr)
            4'b0000 :    data = 16'b00000111_11100000; //
            4'b0001 :    data = 16'b00001111_11110000; //
            4'b0010 :    data = 16'b00001111_11110000; //
            4'b0011 :    data = 16'b00011111_11111000; //
            4'b0100 :    data = 16'b00111111_11111100; //
            4'b0101 :    data = 16'b01111111_11111110; //
            4'b0110 :    data = 16'b11111111_11111111; //
            4'b0111 :    data = 16'b11111111_11111111; //
            4'b1000 :    data = 16'b11111111_11111111; //
            4'b1001 :    data = 16'b11111111_11111111; //
            4'b1010 :    data = 16'b11111111_11111111; //
            4'b1011 :    data = 16'b01111111_11111110; //
            4'b1100 :    data = 16'b00111111_11111100; // 
            4'b1101 :    data = 16'b00011111_11111000; //
            4'b1110 :    data = 16'b00001111_11110000; //
            4'b1111 :    data = 16'b00000111_11100000; // 
        endcase
    
endmodule
